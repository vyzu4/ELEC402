typedef enum logic [2:0] {
    IDLE  = 3'b000,
    WRITE = 3'b001,
    FULL =  3'b010,
    READ = 3'b011,
    EMPTY = 3'b100
} state_t;

module multiplier #(
) (
    input  logic                clk,
    // input  logic                rst,      

    input  logic                EN_mult, // high to start multiplication
    output logic                EN_writeMem, // high to write to mem   
    output logic [6-1:0]        writeMem_addr, // addr to write to

    input  logic [16-1:0]       mult_input0,
    input  logic [16-1:0]       mult_input1,
    output logic [16-1:0]       writeMem_val,  

    output logic                RDY_mult, // ready to multiply             
     
    input  logic                EN_blockRead, // high to read from mem block           
    output logic                VALID_memVal, // high for valid mem val           
    output logic [16-1:0]       memVal_data, // mem data            

    output logic                EN_readMem, // high to start reading mem             
    output logic [6-1:0]        readMem_addr, // addr to read from           
    input  logic [16-1:0]       readMem_val // data read from mem               
);

    state_t state = IDLE;
    state_t next_state;

    // flags
    logic first_write = 1'b0; 
    logic first_read = 1'b0; 
    logic first_VALID_memVal = 1'b0; 

    logic [16-1: 0] product,product_pre;

    // multiplication logic
    always_ff @(posedge clk) begin
        product <= mult_input0 * mult_input1;
        writeMem_val <= product;
    end

    always_comb begin
        memVal_data = readMem_val;   
    end

    // state transition/behaviour logic
    always_ff @(posedge clk) begin
        // next_state = state; // default hold

        // if (!rst)
        //     state = IDLE;
        // else
        //     // transition to next state
        //     state = next_state;

        state = next_state;
        
        unique case (state)

            IDLE: begin
                first_write = 1'b0; //set flag
                
                // initialize write signals
                RDY_mult = 1'b1;
                EN_readMem= 1'b0;
                writeMem_addr = 1'b0;

                // initialize write signals
                readMem_addr = 1'b0;
                VALID_memVal = 1'b0; 

                // determine next state
                if (EN_mult == 1'b1) begin
                    next_state = WRITE;
                end
                else begin
                    next_state = IDLE;
                end
            end

            WRITE: begin
                // initialize write signals
                EN_writeMem = 1'b1;

                // determine value of RDY_mult
                if (writeMem_addr < 6'd61)
                    RDY_mult = 1'b1;
                else
                    RDY_mult = 1'b0;

                // determine EN_writeMem and next state
                if (EN_mult == 1'b0) begin
                    EN_writeMem = 1'b0;
                    next_state = IDLE;
                end
                else begin
                    EN_writeMem = 1'b1;

                    if (writeMem_addr < 6'd62)
                        next_state = WRITE;
                    else
                        next_state = FULL;
                end

                // determine value of writeMem_addr
                writeMem_addr = !first_write ?  1'b0 : writeMem_addr + 1;
                first_write = 1'b1;
            end

            FULL: begin
                // initialize write signals
                RDY_mult = 1'b0;

                first_read = 1'b0; // set flag

                // read related signals
                EN_writeMem = 1'b0;
                writeMem_addr=6'b0;
                EN_readMem = 1'b0;
                readMem_addr = 1'b0;

                // determine next state
                if (EN_mult == 1'b1) begin
                    next_state = FULL;
                end 
                else begin
                    if (EN_blockRead == 1'b1) begin
                        next_state = READ;
                        EN_readMem = 1'b1;
                        readMem_addr = 6'b0;
                    end
                    else 
                        next_state = FULL;
                end
            end

            READ: begin
                // // set flag
                // first_VALID_memVal = 1'b0;

                VALID_memVal = 1'b1;
                // memVal_data <= readMem_val;                
                
                // determine next state
                if (readMem_addr < 6'd63) begin
                    next_state = READ;
                    EN_readMem = 1'b1;
                    readMem_addr =readMem_addr + 1;
                end
                else begin
                    RDY_mult = 1'b1;
                    next_state = IDLE;
                    EN_readMem = 1'b0;
                    // readMem_addr=6'b0;
                end

                // // determine value for VALID_memVal
                // if (EN_readMem == 1'b1)
                //     VALID_memVal = 1'b1;
                // else
                //     VALID_memVal = 1'b0;

                // determine value of writeMem_addr

               //readMem_addr = !first_read ?  1'b0 : readMem_addr + 1;
                // first_read = 1'b1;

            end
/*
            EMPTY: begin
                EN_readMem = 1'b0;
                next_state=IDLE;
                RDY_mult = 1'b1;

                if (EN_mult == 1'b1) 
                    next_state = IDLE;
                else 
                    next_state = EMPTY;

                VALID_memVal = !first_VALID_memVal ?  1'b1 : 1'b0;
                first_VALID_memVal = 1'b1;
            end
            */

            default: next_state = IDLE;
        endcase
    end

endmodule


