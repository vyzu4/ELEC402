`timescale 1ns/1ps
module fsm_tb;
  // multiplier i/o
    logic                clk; // input
    logic                rst; // input     

    logic                EN_mult; // input
    logic                EN_writeMem; // output
    logic [6-1:0]          writeMem_addr; // output

    logic [15:0]         mult_input0; // input
    logic [15:0]         mult_input1; // input
    logic [16-1:0]       writeMem_val; // output 

    logic                RDY_mult;             
     
    logic                EN_blockRead; // input           
    logic                VALID_memVal; // output           
    logic [16-1:0]       memVal_data; // output            

    logic                EN_readMem; // output             
    logic [6-1:0]        readMem_addr; // output           
    logic [16-1:0]       readMem_val; // input 

  /////////////////////////////////////////

    logic           clkA; // input  
    logic           clkB; // input  
    logic [6-1:0]   aA; // input  
    logic [6-1:0]   aB; // input  
    logic           cenA; // input  
    logic           cenB; // input  
    logic [16-1:0]   d; // input  
    logic [16-1:0]   q; // output  

  ////////////////////////////

    // wire            wire_clkA; // input  
    // wire            wire_clkB; // input  
    // wire [6-1:0]    wire_aA; // input  
    // wire [6-1:0]    wire_aB; // input  
    // wire            wire_cenA; // input  
    // wire            wire_cenB; // input  
    // wire [16-1:0]   wire_d; // input  
    // wire [16-1:0]   wire_q; // output  



  // Instantiate multiplier DUT
  multiplier multiplier_dut (
    .clk(clk),
    .rst(rst),

    .EN_mult(EN_mult),
    .EN_writeMem(EN_writeMem),
    .writeMem_addr(writeMem_addr),

    .mult_input0(mult_input0),
    .mult_input1(mult_input1),
    .writeMem_val(writeMem_val),

    .RDY_mult(RDY_mult),

    .EN_blockRead(EN_blockRead),
    .VALID_memVal(VALID_memVal),
    .memVal_data(memVal_data),

    .EN_readMem(EN_readMem),
    .readMem_addr(readMem_addr),
    .readMem_val(q)
  );

  // Instantiate memory_wrapper_2port DUT
  memory_wrapper_2port mw2p_dut (
    .clkA(clk),
    .clkB(clk),

    .aA(readMem_addr),
    .aB(writeMem_addr),

    .cenA(~EN_readMem),
    .cenB(~EN_writeMem),

    .d(writeMem_val),
    .q(q)
  );

  // // Instantiate registerArray DUT
  // registerArray mra_dut (
  //   .clkA(wire_clk),
  //   .clkB(wire_clk),

  //   .aA(wire_readMem_addr),
  //   .aB(wire_writeMem_addr),

  //   .cenA(~wire_EN_readMem),
  //   .cenB(~wire_EN_writeMem),

  //   .d(wire_writeMem_val),
  //   .q(wire_q)
  // );


  // Clock generator
  initial clk = 0;
  always #1.25 clk = ~clk; // 400 MHz
  // always #0.625 clk = ~clk; // 800 MHz

  always begin
    #10 mult_input0 = 16'd1; mult_input1 = 16'd9;
    #10 mult_input0 = 16'd2; mult_input1 = 16'd8;
    #10 mult_input0 = 16'd3; mult_input1 = 16'd7;
    #10 mult_input0 = 16'd4; mult_input1 = 16'd6;
    #10 mult_input0 = 16'd5; mult_input1 = 16'd5;
    #10 mult_input0 = 16'd6; mult_input1 = 16'd4;
    #10 mult_input0 = 16'd7; mult_input1 = 16'd3;
    #10 mult_input0 = 16'd8; mult_input1 = 16'd2;
    #10 mult_input0 = 16'd9; mult_input1 = 16'd1;
  end

  // Stimulus to fsm
  initial begin
    // initialize signals
    #10 rst = 1; EN_mult = 0; EN_blockRead = 0; 
    #10 rst = 0;
    #10 EN_mult = 1;            
    #700;
    #10 EN_mult = 0; // stop writing
    #10 EN_blockRead = 1;
    #10 EN_blockRead = 0;

    #700 EN_mult = 1;
    #700;

    $stop;
  end

endmodule

